module clock;