module timing