module counting;